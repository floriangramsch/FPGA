--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ex03_lfsr8_tb is
generic (
    g_CLK_MHZ : real := 1000.0--;
);
end entity;

architecture arch of ex03_lfsr8_tb is

    signal clk : std_logic := '1';
    signal reset_n : std_logic := '0';
    signal cycle : integer := 0;

    -- define constant array C_LFSR8_SEQUENCE of 256 8-bit vectors
    -- and initialize it with the sequence provided in lfsr8.txt
    type array_8b_t is array (natural range <>) of std_logic_vector(7 downto 0);
    constant C_LFSR8_SEQUENCE : array_8b_t(0 to 255) := (
        "00000000",        "00000001",        "00000011",        "00000111",        "00001111",        "00011110",        "00111101",        "01111010",
        "11110100",        "11101000",        "11010000",        "10100001",        "01000011",        "10000111",        "00001110",        "00011100",
        "00111001",        "01110010",        "11100101",        "11001011",        "10010111",        "00101111",        "01011111",        "10111111",
        "01111111",        "11111110",        "11111101",        "11111011",        "11110111",        "11101110",        "11011100",        "10111000",
        "01110001",        "11100011",        "11000111",        "10001110",        "00011101",        "00111011",        "01110110",        "11101101",
        "11011010",        "10110100",        "01101000",        "11010001",        "10100011",        "01000111",        "10001111",        "00011111",
        "00111111",        "01111110",        "11111100",        "11111001",        "11110011",        "11100110",        "11001101",        "10011011",
        "00110110",        "01101101",        "11011011",        "10110110",        "01101100",        "11011001",        "10110010",        "01100100",
        "11001000",        "10010001",        "00100011",        "01000110",        "10001101",        "00011011",        "00110111",        "01101111",
        "11011111",        "10111110",        "01111101",        "11111010",        "11110101",        "11101010",        "11010100",        "10101001",
        "01010010",        "10100100",        "01001001",        "10010010",        "00100101",        "01001010",        "10010100",        "00101001",
        "01010011",        "10100110",        "01001101",        "10011010",        "00110100",        "01101001",        "11010011",        "10100111",
        "01001111",        "10011110",        "00111100",        "01111000",        "11110000",        "11100000",        "11000001",        "10000010",
        "00000100",        "00001001",        "00010010",        "00100100",        "01001000",        "10010000",        "00100001",        "01000010",
        "10000101",        "00001010",        "00010100",        "00101000",        "01010001",        "10100010",        "01000101",        "10001011",
        "00010111",        "00101110",        "01011101",        "10111011",        "01110111",        "11101111",        "11011110",        "10111100",
        "01111001",        "11110010",        "11100100",        "11001001",        "10010011",        "00100111",        "01001110",        "10011100",
        "00111000",        "01110000",        "11100001",        "11000011",        "10000110",        "00001100",        "00011000",        "00110001",
        "01100011",        "11000110",        "10001100",        "00011001",        "00110011",        "01100111",        "11001110",        "10011101",
        "00111010",        "01110100",        "11101001",        "11010010",        "10100101",        "01001011",        "10010110",        "00101101",
        "01011011",        "10110111",        "01101110",        "11011101",        "10111010",        "01110101",        "11101011",        "11010110",
        "10101101",        "01011010",        "10110101",        "01101010",        "11010101",        "10101011",        "01010110",        "10101100",
        "01011000",        "10110001",        "01100010",        "11000100",        "10001000",        "00010001",        "00100010",        "01000100",
        "10001001",        "00010011",        "00100110",        "01001100",        "10011000",        "00110000",        "01100001",        "11000010",
        "10000100",        "00001000",        "00010000",        "00100000",        "01000000",        "10000001",        "00000010",        "00000101",
        "00001011",        "00010110",        "00101100",        "01011001",        "10110011",        "01100110",        "11001100",        "10011001",
        "00110010",        "01100101",        "11001010",        "10010101",        "00101011",        "01010111",        "10101110",        "01011100",
        "10111001",        "01110011",        "11100111",        "11001111",        "10011111",        "00111110",        "01111100",        "11111000",
        "11110001",        "11100010",        "11000101",        "10001010",        "00010101",        "00101010",        "01010101",        "10101010",
        "01010100",        "10101000",        "01010000",        "10100000",        "01000001",        "10000011",        "00000110",        "00001101",
        "00011010",        "00110101",        "01101011",        "11010111",        "10101111",        "01011110",        "10111101",        "01111011",
        "11110110",        "11101100",        "11011000",        "10110000",        "01100000",        "11000000",        "10000000",        "00000000"
    );

    signal s_sequence_cntr : integer := 0;

    -- create an array of 256 unsigned integers (natural)
    -- and initialize all elements to zero
    type array_natural_t is array (natural range <>) of natural;
     -- this array will store the number of times the lfsr value was seen
    signal s_lfsr_value : array_natural_t(0 to 255) := (others => 0);

    signal lfsr, period : std_logic_vector(7 downto 0);

begin

    clk <= not clk after (0.5 us / g_CLK_MHZ);
    reset_n <= '0', '1' after (2.0 us / g_CLK_MHZ);
    cycle <= cycle + 1 after (1 us / g_CLK_MHZ);

    e_lfsr8 : entity work.ex03_lfsr8
    port map (
        o_lfsr => lfsr,
        o_period => period,
        i_reset_n => reset_n,
        i_clk => clk--,
    );

    process(clk, reset_n)
    begin
    if ( reset_n = '0' ) then
        --
    elsif rising_edge(clk) then
        -- in the simulation check, look-up the expected value in the constant array (based on the current position in the sequence)
        -- and stop the simulation when there is a mismatch
        assert ( lfsr = C_LFSR8_SEQUENCE(s_sequence_cntr mod 255) ) severity error;

        -- increment a counter s_sequence_cntr to count the current position in the sequence
        s_sequence_cntr <= s_sequence_cntr + 1;

        -- increment s_lfsr_value's element of the current LFSR value to count how often a value appears during a sequence
        s_lfsr_value(to_integer(unsigned(lfsr))) <= s_lfsr_value(to_integer(unsigned(lfsr))) + 1;

        if ( s_sequence_cntr = 255 ) then
            report "Simulation DONE";
        end if;
        --
    end if;
    end process;

end architecture;
